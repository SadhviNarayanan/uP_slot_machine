module rom_wrapper (
    input  logic clk,
    input  logic [2:0] sprite_idx,       // 0-6 for 7 sprites
    input  logic [5:0] x_in_sprite,      // 0-63
    input  logic [5:0] y_in_sprite,      // 0-63
    output logic [2:0] pixel_rgb         // 3-bit RGB output
);

    localparam SPRITE_WIDTH = 64;
    localparam SPRITE_HEIGHT = 64;

    // 28 BRAMs total (4 per sprite × 7 sprites)
    // Each word stores 5 pixels (5 × 3 = 15 bits, 1 bit unused)
    logic [15:0] bram [0:27][0:255]; // 256x16 BRAMS -- 256 lines, 16bit words
    
    // Load sprite data
    initial begin
        $readmemh("sprite0_bram0.mem", bram[0]);
        $readmemh("sprite0_bram1.mem", bram[1]);
        $readmemh("sprite0_bram2.mem", bram[2]);
        $readmemh("sprite0_bram3.mem", bram[3]);
        
        $readmemh("sprite1_bram0.mem", bram[4]);
        $readmemh("sprite1_bram1.mem", bram[5]);
        $readmemh("sprite1_bram2.mem", bram[6]);
        $readmemh("sprite1_bram3.mem", bram[7]);
        
        $readmemh("sprite2_bram0.mem", bram[8]);
        $readmemh("sprite2_bram1.mem", bram[9]);
        $readmemh("sprite2_bram2.mem", bram[10]);
        $readmemh("sprite2_bram3.mem", bram[11]);
        
        $readmemh("sprite3_bram0.mem", bram[12]);
        $readmemh("sprite3_bram1.mem", bram[13]);
        $readmemh("sprite3_bram2.mem", bram[14]);
        $readmemh("sprite3_bram3.mem", bram[15]);
        
        $readmemh("sprite4_bram0.mem", bram[16]);
        $readmemh("sprite4_bram1.mem", bram[17]);
        $readmemh("sprite4_bram2.mem", bram[18]);
        $readmemh("sprite4_bram3.mem", bram[19]);
        
        $readmemh("sprite5_bram0.mem", bram[20]);
        $readmemh("sprite5_bram1.mem", bram[21]);
        $readmemh("sprite5_bram2.mem", bram[22]);
        $readmemh("sprite5_bram3.mem", bram[23]);
        
        $readmemh("sprite6_bram0.mem", bram[24]);
        $readmemh("sprite6_bram1.mem", bram[25]);
        $readmemh("sprite6_bram2.mem", bram[26]);
        $readmemh("sprite6_bram3.mem", bram[27]);
    end
    
    // Calculate pixel index within sprite (0-4095)
    // NOTE: this is just for pixels of which there are 4096 - each of these have 3 bits for rgb which are stored in memory hence we need 4
    // so when are doing calcualtions we want to treat it as pixels and not bits - hence we abstract away each bit (treat as 5 insted of 5*3=15 for example)
    logic [11:0] pixel_index;
    assign pixel_index = (y_in_sprite * SPRITE_WIDTH) + x_in_sprite;
    // Example: y=2, x=25 → pixel_index = 2*64 + 25 = 153
    
    // Divide by 5 to get word offset within sprite -- which word line??
    logic [11:0] word_offset;
    assign word_offset = pixel_index / 5;
    
    // Which of the 4 BRAMs for this sprite? --> got which word line its own, now need to see which block this wordline belowngs to
    logic [1:0] bram_offset;    // 0-3
    assign bram_offset = word_offset[9:8];  // word_offset / 256 --> essetnailly dividing pixel_index / (# of pixels in a block), where # of pixels in a block is number of words * 5 = 256 * 5 (since 5 pixels in a word line)
    
    // Address within that BRAM
    logic [7:0] bram_addr;
    assign bram_addr = word_offset[7:0];    // word_offset % 256 --> remainder of the division above, essentiallu tells us spill over into RAM block since it doesn't alsways divide eprfectly into a block   

    // Absolute BRAM index (0-27)
    logic [4:0] bram_index;
    assign bram_index = (sprite_idx << 2) + bram_offset;  // sprite_idx * 4 + bram_offset --> since each index gets 4 blocks
    
    // Which of 5 pixels in the word?
    logic [2:0] pixel_in_word;
    assign pixel_in_word = pixel_index % 5;


    
    logic [15:0] selected_word;
    
    always_ff @(posedge clk) begin
        // Read from the calculated BRAM and address
        selected_word <= bram[bram_index][bram_addr];
        
        // Extract the right 3-bit pixel from the word
        // Word format: [15]=unused, [14:12]=pix4, [11:9]=pix3, [8:6]=pix2, [5:3]=pix1, [2:0]=pix0
        case (pixel_in_word)
            3'd0: pixel_rgb <= selected_word[2:0];
            3'd1: pixel_rgb <= selected_word[5:3];
            3'd2: pixel_rgb <= selected_word[8:6];
            3'd3: pixel_rgb <= selected_word[11:9]; 
            3'd4: pixel_rgb <= selected_word[14:12];
            default: pixel_rgb <= 3'b000;
        endcase
    end

endmodule